module Controller_Cancela( Cancela, GO);
  input GO;
  output Cancela;
  
  assign Cancela = GO;
 
endmodule 